library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity MEMORIA_PROGRAMA00 is
    Port ( A : in  STD_LOGIC_VECTOR (5 downto 0);
           D : out  STD_LOGIC_VECTOR (31 downto 0));
end MEMORIA_PROGRAMA00;

architecture MEMORIA_PROGRAMA0 of MEMORIA_PROGRAMA00 is

-- CARGA Y ALMACENAMIENTO
	CONSTANT OPCODE_LW	 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000";
	CONSTANT OPCODE_SW		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00001";

-- OPERACIONES ARITMETICAS
	CONSTANT OPCODE_SUM 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00010";
	CONSTANT OPCODE_REST 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00011";
	CONSTANT OPCODE_MULT 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00100";
	
--OPERACIONES LOGICAS
	CONSTANT OPCODE_AND 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00101";
	CONSTANT OPCODE_OR   	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00110";
	CONSTANT OPCODE_NOT 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00111";
	CONSTANT OPCODE_XOR 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01000";
	CONSTANT OPCODE_XNOR 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01001";
	CONSTANT OPCODE_NAND 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01010";
	CONSTANT OPCODE_NOR 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01011";
	
--OPERACIONES COMPARADOR
	CONSTANT OPCODE_MYQ 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01100";
	CONSTANT OPCODE_MNQ 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01101";
	CONSTANT OPCODE_IGU 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01110";
	CONSTANT OPCODE_MYI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01111";
	CONSTANT OPCODE_MNI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10001";
	CONSTANT OPCODE_DIF 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10010";
	
-- SALTOS	
	CONSTANT OPCODE_B	 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10011";
	CONSTANT OPCODE_BNEQ	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10100";

-- REGISTROS	
	CONSTANT R0					: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	CONSTANT R1					: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000001";
	CONSTANT R2					: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000010";
	CONSTANT R3					: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000011";
	CONSTANT R4					: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000100";
	CONSTANT R5					: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000101";
	CONSTANT R6					: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000110";
	CONSTANT R7					: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000111";
	CONSTANT R8					: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00001000";
	CONSTANT R9					: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00001001";
	CONSTANT R10				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00001010";
	CONSTANT R11				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00001011";
	CONSTANT R12				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00001100";
	CONSTANT R13				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00001101";
	CONSTANT R14				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00001110";
	CONSTANT R15				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00001111";
	CONSTANT R16				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00010000";
	CONSTANT R17				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00010001";
	CONSTANT R18				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00010010";
	CONSTANT R19				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00010011";
	CONSTANT R20				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00010100";
	CONSTANT R21				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00010101";
	CONSTANT R22				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00010110";
	CONSTANT R23				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00010111";
	CONSTANT R24				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00011000";
	CONSTANT R25				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00011001";
	CONSTANT R26				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00011010";
	CONSTANT R27				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00011011";
	CONSTANT R28				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00011100";
	CONSTANT R29				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00011101";
	CONSTANT R30				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00011110";
	CONSTANT R31				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00011111";
	CONSTANT R32				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00100000";
	CONSTANT R33				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00100001";
	CONSTANT R34				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00100010";
	CONSTANT R35				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00100011";
	CONSTANT R36				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00100100";
	CONSTANT R37				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00100101";
	CONSTANT R38				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00100110";
	CONSTANT R39				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00100111";
	CONSTANT R40				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00101000";
	CONSTANT R41				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00101001";
	CONSTANT R42				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00101010";
	CONSTANT R43				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00101011";
	CONSTANT R44				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00101100";
	CONSTANT R45				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00101101";
	CONSTANT R46				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00101110";
	CONSTANT R47				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00101111";
	CONSTANT R48				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00110000";
	CONSTANT R49				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00110001";
	CONSTANT R50				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00110010";
	CONSTANT R51				: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00110011";

-- SIN USO
	CONSTANT SU					: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	
-- INICIO DIRECCION 	
	CONSTANT CR				: STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";	

	
	TYPE ARR IS ARRAY (0 TO 256) OF STD_LOGIC_VECTOR(31 DOWNTO 0); 
	CONSTANT ROM : ARR := (
	
	OPCODE_LW & R0 & SU & "00000000101",	 	
	OPCODE_SW & SU & R1 & "00000000110", 
	
	OPCODE_SUM & R2 & R3 & R4 & CR, 
	OPCODE_REST & R5 & R6 & R7 & CR,	
	OPCODE_MULT & R8 & R9 & R10 & CR,	
	OPCODE_AND & R11 & R12 & R13 & CR,
	OPCODE_OR & R14 & R15 & R16 & CR,  	
	OPCODE_NOT & R17 & R18 & R19 & CR,	
	OPCODE_XOR & R20 & R21 & R22 & CR,	
	OPCODE_XNOR & R23 & R24 & R25 & CR,	
	OPCODE_NAND & R26 & R27 & R28 & CR,	
	OPCODE_NOR & R29 & R30 & R31 & CR,	
	OPCODE_MYQ & R32 & R33 & R34 & CR,	
	OPCODE_MNQ & R35 & R36 & R37 & CR,	
	OPCODE_IGU & R38 & R39 & R40 & CR,	
	OPCODE_MYI & R41 & R42 & R43 & CR,
	OPCODE_MNI & R44 & R45 & R46 & CR,	
	OPCODE_DIF & R47 & R48 & R49 & CR,
	
	OPCODE_BNEQ	& R50 & R51 &"00000001000",
	OPCODE_B & SU & SU & "00000000111",	
	
	
		
		OTHERS=>(OTHERS=>'0')
	);
begin
	D <= ROM( CONV_INTEGER(A) );
end MEMORIA_PROGRAMA0;

